library ieee;
use ieee.std_logic_1164.all;

package sim_aurora_pkg is
	type tData is array(natural range <>) of std_logic_vector(7 downto 0);
end package;
